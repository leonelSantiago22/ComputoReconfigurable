//unidad de control
module fetch #(parameter N=3)
(
		input logic [3*N+2:0]dout,
		output logic [N-1:0] d0,d1,
		output logic [2:0] a0,a1
		output logic we
);

	always_comb
			
endmodule
