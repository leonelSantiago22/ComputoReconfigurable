module practica1(input logic 
